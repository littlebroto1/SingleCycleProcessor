../../../ControlUnit/hdl/sv/Decoder.sv