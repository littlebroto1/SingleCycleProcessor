../../../Mux2/hdl/sv/mux2.sv