../../../Extender/hdl/sv/extender.sv