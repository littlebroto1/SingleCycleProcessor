../../../ControlUnit/hdl/sv/MainDecoder.sv