../../../RAM/hdl/sv/ram.sv