../../../PCLogic/hdl/sv/PCLogic.sv