../../../Shift/hdl/sv/shift.sv