../../../ConditionLogic/hdl/sv/ConditionLogic.sv