../../../Decoder/hdl/sv/Decoder.sv