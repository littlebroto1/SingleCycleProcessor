../../../ControlUnit/hdl/sv/EnabledFF.sv