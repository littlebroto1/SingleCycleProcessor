../../../ConditionCheck/hdl/sv/ConditionCheck.sv