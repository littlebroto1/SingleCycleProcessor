../../../ALU/hdl/sv/alu.sv