../../../ALUDecoder/hdl/sv/ALUDecoder.sv