../../../MainDecoder/hdl/sv/MainDecoder.sv