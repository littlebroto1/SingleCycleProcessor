../../../ControlUnit/hdl/sv/PCLogic.sv