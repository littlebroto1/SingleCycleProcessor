../../../ControlUnit/hdl/sv/ConditionCheck.sv