../../../RegisterFile/hdl/sv/registerfile.sv