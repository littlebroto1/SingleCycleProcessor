../../../ControlUnit/hdl/sv/ControlUnit.sv