../../../EnabledFF/hdl/sv/EnabledFF.sv