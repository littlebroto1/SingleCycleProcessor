../../../ControlUnit/hdl/sv/ConditionLogic.sv