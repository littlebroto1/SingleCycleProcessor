../../../ControlUnit/hdl/sv/ALUDecoder.sv